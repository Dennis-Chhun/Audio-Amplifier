**************************************
.end
