
* LM317MOT Voltage Reg. (Motorola)
*
.SUBCKT LM317MOT 1      2    3
*Connections  Input  Adj. Output
*LM317A voltage regulator - Motorola
J1 1 3 4 JN
Q2 5 5 6 QPL .1
Q3 5 8 9 QNL  .2
Q4 8 5 7 QPL .1
Q5 81 8 3 QNL .2
Q6 3 81 10 QPL .2
Q7 12 81 13 QNL  .2
Q8 10 5 11 QPL  .2
Q9 14 12 10 QPL .2
Q10 16 5 17 QPL  .2
Q11 16 14 15 QNL .2
Q12 3 20 16 QPL .2
Q13 1 19 20 QNL .2
Q14 19 5 18 QPL .2
Q15 3 21 19 QPL .2
Q16 21 22 16 QPL .2
Q17 21 3 24 QNL   .2
Q18 22 22 16 QPL .2
Q19 22 3 241 QNL 2
Q20 3 25 16 QPL .2
Q21 25 26 3 QNL .2
Q22A 35 35 1 QPL 2
Q22B 16 35 1 QPL 2
Q23 35 16 30 QNL  2
Q24A 27 40 29 QNL .2
Q24B 27 40 28 QNL .2
Q25 1 31 41 QNL 5
Q26 1 41 32 QNL 50
D1 3 4 DZ
D2 33 1 DZ
D3 29 34 DZ
R1 1 6 310
R2 1 7 310
R3 1 11 230
R4 1 17 120
R5 1 18 5.6K
R6 4 8 125K
R7 8 81 135
R8 10 12 12.4K
R9 9 3 190
R10 13 3 3.6K
R11 14 3 5.8K
R12 15 3 110
R13 20 3 5.1K
R14 2 24 12.5K
R15 24 241 2.4K
R16 16 25 6.7K
R17 16 40 12K
R18 30 41 160
R19 16 31 170
R20 26 27 6.8K
R21 27 40 510
R22 3 41 200
R23 33 34 13K
R24 28 29 105
R25 28 32 4
R26 32 3 .1
C1 21 3 30PF
C2 21 2 30PF
C3 25 26 5PF
CBS1 5 3 2PF
CBS2 35 3 1PF
CBS3 22 3 1PF
.MODEL JN NJF(BETA=1E-4 VTO=-7)
.MODEL DZ D(BV=6.3)
.MODEL QNL NPN(EG=1.22 BF=80 RB=100 CCS=1.5PF TF=.3NS TR=6NS CJE=2PF
+ CJC=1PF VAF=100)
.MODEL QPL PNP(BF=40 RB=20 TF=.6NS TR=10NS CJE=1.5PF CJC=1PF VAF=50)
.ENDS LM317MOT
*
